//###########################################################################
//
//  Copyright 2021 The SVUnit Authors.
//
//  Licensed under the Apache License, Version 2.0 (the "License");
//  you may not use this file except in compliance with the License.
//  You may obtain a copy of the License at
//
//      http://www.apache.org/licenses/LICENSE-2.0
//
//  Unless required by applicable law or agreed to in writing, software
//  distributed under the License is distributed on an "AS IS" BASIS,
//  WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
//  See the License for the specific language governing permissions and
//  limitations under the License.
//
//###########################################################################

package junit_xml;

  `include "XmlElement.svh"
  `include "TestCase.svh"
  `include "TestSuite.svh"

  // test_suites[] needs to be declared as a dynamic array[$] (not a static array[] with a fixed length)
  //
  function automatic string to_xml_report_string(input TestSuite test_suites[$]);
    XmlElement testsuites = new("testsuites");
    foreach (test_suites[i])
      testsuites.add_child(test_suites[i].as_xml_element());
    return testsuites.as_string();
  endfunction

endpackage
